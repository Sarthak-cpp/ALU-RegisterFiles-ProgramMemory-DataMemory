LIBRARY IEEE;
    USE IEEE.STD_LOGIC_1164.ALL;
    USE IEEE.STD_LOGIC_UNSIGNED.ALL;
    USE IEEE.NUMERIC_STD.ALL;

--Program Memory Design
Entity ProgramMemory IS
	PORT(
    	add: IN STD_LOGIC_VECTOR(5 downto 0);
        RDat: OUT STD_LOGIC_VECTOR(31 downto 0)
        );
End Entity;

--Program Memory Architecture

Architecture BEV of ProgramMemory IS
TYPE MEM IS ARRAY (63 DOWNTO 0) OF STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL MEMORY : MEM:=("11000010101110001001101000111010",
"01001110011100011101001010110000",
"00100101111010000110101010100100",
"10111011101000011001001001000011",
"00011110000101001101001000001001",
"10101010111110111011000110010011",
"11000110001110110011100010001101",
"11111001101101001011010100101110",
"11100000001001011111111111101001",
"11111010100011111101010110111110",
"01101000000100100000011010110010",
"10101001011001100000010110010010",
"00110001011110100010111110010000",
"00100000000001010001010110010011",
"00000111101111111110011010010001",
"00000101000111000111011111010010",
"11010010101110010010100101111101",
"11000111101110111111110001000011",
"11111110001011010101000111001011",
"00000100110001100011110110111101",
"01001011111000011001010011100101",
"11110101101101010011011010000000",
"01101110000010011111100101010101",
"01110011111110111100001001011110",
"11101111011100001000011110011011",
"00101111010001110101111101110001",
"10001100100011100000000001010000",
"01000000001110111010010010100001",
"00010011100111010000111000111011",
"01001011001000110000111000011001",
"01100011000011111111000011110001",
"11010000101001101010111000010111",
"11100011011100011101110001100010",
"00010101111100111000110110101001",
"10110111010010000000111001000100",
"01101001000001111100101100010000",
"11000010011111110100110011100011",
"11011000001101011000110000101110",
"00011100011001101010011001111000",
"11010011100010001110111001110011",
"10001101110011010000001010011001",
"00011101011101100000111000001011",
"11000010101001011111101010000001",
"10001011011010001001110010010111",
"00101011011111110000101011011001",
"11011001011110011010101100100010",
"01110010100101000001110100011110",
"10000101010111110101110100111100",
"11110110001111111101111111100011",
"01011001001100100101110011000010",
"00110000000010100110010101011100",
"10111000100010100001001100110110",
"01111100111100011110001000100011",
"01101011110100001100100011100110",
"00110010110011001100101001001000",
"10001001010110001010111111001101",
"00100010110000101001110101011111",
"01110100010110111010000101000111",
"11111001010111111111010110011101",
"10001001101010100010101110100101",
"01010111110000111011001110111110",
"00011111100100010000110010010110",
"11000000010101110101011000100100",
"10100001001000011001000100101001")
;
SIGNAL ADDR : INTEGER RANGE 0 TO 63;

Begin
	Process(add)
    Begin
    ADDR<=CONV_INTEGER(add);
    RDat<=MEMORY(ADDR);
    End Process;
End BEV;